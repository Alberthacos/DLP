----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:21:13 09/04/2022 
-- Design Name: 
-- Module Name:    d - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity d is
    Port ( a : in  STD_LOGIC;
           AS : in  STD_LOGIC;
           D : in  STD_LOGIC;
           S : in  STD_LOGIC;
           D : in  STD_LOGIC_VECTOR (3 downto 1);
           A : in  STD_LOGIC);
end d;

architecture Behavioral of d is

begin


end Behavioral;

